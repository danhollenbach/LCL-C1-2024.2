module starter(
input clk,
output data
);

endmodule