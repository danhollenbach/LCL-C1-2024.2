library verilog;
use verilog.vl_types.all;
entity Pre3_vlg_vec_tst is
end Pre3_vlg_vec_tst;
