module zeroer(
output [6:0] out
);

// designa a saida dos displays de 7 segmentos nao usados para 1 e os apaga
assign out = 7'b1111111;

endmodule
