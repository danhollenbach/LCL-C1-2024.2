library verilog;
use verilog.vl_types.all;
entity Exp52_vlg_vec_tst is
end Exp52_vlg_vec_tst;
