library verilog;
use verilog.vl_types.all;
entity Pre2 is
    port(
        B0              : out    vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        B1              : out    vl_logic;
        B3              : out    vl_logic;
        B4              : out    vl_logic;
        B5              : out    vl_logic;
        B6              : out    vl_logic;
        B7              : out    vl_logic;
        B8              : out    vl_logic;
        B9              : out    vl_logic;
        B2              : out    vl_logic
    );
end Pre2;
