library verilog;
use verilog.vl_types.all;
entity Exp53_vlg_vec_tst is
end Exp53_vlg_vec_tst;
