library verilog;
use verilog.vl_types.all;
entity Exp53_vlg_check_tst is
    port(
        S               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Exp53_vlg_check_tst;
