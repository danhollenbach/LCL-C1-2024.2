library verilog;
use verilog.vl_types.all;
entity Exp51_vlg_check_tst is
    port(
        COUT            : in     vl_logic;
        SUM             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Exp51_vlg_check_tst;
