library verilog;
use verilog.vl_types.all;
entity exp8_vlg_check_tst is
    port(
        COUNT           : in     vl_logic_vector(2 downto 0);
        sampler_rx      : in     vl_logic
    );
end exp8_vlg_check_tst;
