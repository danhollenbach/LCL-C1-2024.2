library verilog;
use verilog.vl_types.all;
entity Exp10_vlg_vec_tst is
end Exp10_vlg_vec_tst;
