module opcreator(
input clk, 
input [2:0] op,
output [2:0] result
);

always_ff @(posedge clk)
result <= op;

endmodule 