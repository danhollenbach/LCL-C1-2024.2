library verilog;
use verilog.vl_types.all;
entity Pre2_vlg_vec_tst is
end Pre2_vlg_vec_tst;
