module senha (
output [6:0] seed
);

assign seed = 7'b1101101;

endmodule