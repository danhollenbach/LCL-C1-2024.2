library verilog;
use verilog.vl_types.all;
entity Exp51_vlg_vec_tst is
end Exp51_vlg_vec_tst;
