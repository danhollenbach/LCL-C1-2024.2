library verilog;
use verilog.vl_types.all;
entity Pre1_vlg_vec_tst is
end Pre1_vlg_vec_tst;
