library verilog;
use verilog.vl_types.all;
entity Pre2_vlg_check_tst is
    port(
        B0              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        B3              : in     vl_logic;
        B4              : in     vl_logic;
        B5              : in     vl_logic;
        B6              : in     vl_logic;
        B7              : in     vl_logic;
        B8              : in     vl_logic;
        B9              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Pre2_vlg_check_tst;
