module zeroer(
output [6:0] out
);

assign out = 7'b1111111;

endmodule
